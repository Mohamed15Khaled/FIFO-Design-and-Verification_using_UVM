package shared_pkg ;
    int error_count  ;
    int correct_count  ; 
    logic test_finished ;
endpackage